** Profile: "SCHEMATIC1-time_domain"  [ D:\SPB_DATA\APII_LAB3\apii_lab3-pspicefiles\schematic1\time_domain.sim ] 

** Creating circuit file "time_domain.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "D:/Cadence/SPB_16.5/tools/pspice/library/ebipolar.lib" 
* From [PSPICE NETLIST] section of D:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
